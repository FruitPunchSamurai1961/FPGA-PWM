-- PWM_GEN.VHD (a peripheral module for SCOMP)
-- 2021.03.20
--
-- Generates a square wave with duty cycle dependant on value
-- sent from SCOMP.

LIBRARY IEEE;
LIBRARY LPM;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE LPM.LPM_COMPONENTS.ALL;

ENTITY PWM_GEN IS
    PORT(PWMCLOCK,
        RESETN,
        CS       : IN STD_LOGIC;
        IO_DATA  : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		  IN1		  : OUT STD_LOGIC;
		  IN2      : OUT STD_LOGIC;
		  STBY	  : OUT STD_LOGIC;
        PWM_OUT  : OUT STD_LOGIC;
		  IO_WRITE    : IN    STD_LOGIC

    );
END PWM_GEN;

ARCHITECTURE a OF PWM_GEN IS
    SIGNAL COUNT    : STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL COMPARE  : STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL AB	     : STD_LOGIC_VECTOR(1 downto 0);
	 SIGNAL PWM		  : STD_LOGIC;
	 
	
	BEGIN
    IO_Handler: PROCESS (RESETN, CS,IO_WRITE,IO_DATA)
    BEGIN
        -- Create a register to store the data sent from SCOMP
        IF (RESETN = '0') THEN
            COMPARE <= "0000";
				AB <= "00";
        ELSIF (rising_edge(CS) AND IO_WRITE = '1') THEN
            -- When written to, latch IO_DATA into the compare register.
            COMPARE <= IO_DATA(3 DOWNTO 0);
				AB <= IO_DATA(5 DOWNTO 4);
        END IF;

    END PROCESS;

    PWM_Generator: PROCESS (RESETN, PWMCLOCK)
    BEGIN
        -- Something to consider (eventually): should anything happen at reset?
		  IF (RESETN = '0') THEN
				COUNT <= "0000";
				PWM <= '1';
        -- Create a counter and a comparator that control the output
        ELSIF (rising_edge(PWMCLOCK)) THEN
				COUNT <= COUNT + 1;
            -- todo: on compare match, set the output low.
				IF COMPARE = "1111" THEN
					PWM <= '1';
				ELSIF COMPARE = "0000" THEN
					PWM <= '0';
				ELSIF COUNT = COMPARE THEN
					PWM <= '0';
				ELSIF COUNT = "0000" THEN
					PWM <= '1';
				END IF;
        END IF;
    END PROCESS;
	PWM_OUT <= PWM;
	IN1 <= AB(1);
	IN2 <= AB(0);
	STBY <= '0' WHEN (RESETN = '0' OR (AB(0) = '0' AND AB(1) = '0')) ELSE '1';
END a;